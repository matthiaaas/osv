module main

@[export: "kmain"]
fn kmain() {
	for {}
}
