// module main

// pub enum ProcState {
// 	unused
// 	running
// 	sleeping
// 	zombie
// }

// pub struct Process {
// 	pid u32
// 	state ProcState
// 	pagetable Pagetable
// 	kernel_sp voidptr
// }

// pub fn Process.new(pid u32, stack_top voidptr) Process {
// 	return Process{
// 		pid: pid
// 		state: .ready
// 		stack_top: stack_top
// 	}
// }
