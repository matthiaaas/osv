module proc

pub struct Dispatcher {
}

pub fn (mut dispatcher Dispatcher) run(process Process) {
}
