module main

pub struct String {
}

pub fn String.empty() String {
	return String{}
}

pub fn (s String) next() ?u8 {
	return 72
}
