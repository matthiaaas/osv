module memory

pub struct Pagetable {}
