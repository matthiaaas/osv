module trap

@[export: "trap_handler"]
fn trap_handler() {
	for {}
}
