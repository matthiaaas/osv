module proc

pub struct Scheduler {
mut:
	processes [64]Process
}
